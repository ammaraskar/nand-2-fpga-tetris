module not_1(output wire Y, input wire A);
    nand_2 inverter(Y, A, A);
endmodule
